* C:\Users\Theje\eSim-Workspace\Clock_Gating_with_Muller_C\Clock_Gating_with_Muller_C.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/23/26 18:08:07

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ muller_c		
U6  Net-_U3-Pad3_ Net-_U6-Pad2_ Net-_U6-Pad3_ muller_c		
U7  Net-_U4-Pad3_ Net-_U6-Pad2_ d_buffer		
U5  Net-_U4-Pad3_ Net-_U3-Pad1_ d_inverter		
v1  clk GND pulse		
v2  en GND pulse		
U9  Net-_U6-Pad3_ Net-_U8-Pad2_ Net-_U10-Pad1_ d_and		
U8  Net-_U6-Pad2_ Net-_U8-Pad2_ d_buffer		
U4  clk en Net-_U4-Pad3_ Net-_U3-Pad2_ adc_bridge_2		
U10  Net-_U10-Pad1_ clkg dac_bridge_1		
U1  clk plot_v1		
U2  en plot_v1		
U11  clkg plot_v1		

.end
